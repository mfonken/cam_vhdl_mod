library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package global_constants is

-- Ora defaults
	constant DEFAULT_THRESH : integer 	:= 200;
	constant DEFAULT_KERNEL : integer 	:= 0;


end global_constants;
