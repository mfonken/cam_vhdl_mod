library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.ora_types.all;

package ora_constants is


end ora_constants;
