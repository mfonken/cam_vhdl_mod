library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package global_constants is

-- Camera info
	constant OV9712_ADDR : std_logic_vector( 6 downto 0 ) := b"0000000"; -- TODO: get actual address
	


end global_constants;